//----------------------+-------------------------------------------------------
// Filename             | uart_ctrl.vh
// File created on      | 14/06/2022 12:48:12
// Created by           | Sree Sankar E
//                      |
//                      |
//                      |
//----------------------+-------------------------------------------------------
//
//------------------------------------------------------------------------------
// Header of UART Controller
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Register Offset Map
//------------------------------------------------------------------------------

`define CTRL_REG_ADDR       32'h0000_0000
`define STATUS_REG_ADDR     32'h0000_0004
`define TX_DATA_REG_ADDR    32'h0000_0008
`define RX_DATA_REG_ADDR    32'h0000_000C