//----------------------+-------------------------------------------------------
// Filename             | memory_map.vh
// File created on      | 15.11.2020 12:07:34
// Created by           | Sree Sankar E
//                      |
//                      |
//                      |
//----------------------+-------------------------------------------------------
//
//------------------------------------------------------------------------------
// Memory Map
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// OCM
//------------------------------------------------------------------------------

`define OCM_BASE_ADDR       32'h0000_0000
`define OCM_OFFSET          32'h0000_FFFF

//------------------------------------------------------------------------------
// Pheripherals
//------------------------------------------------------------------------------

// UART 0
`define UART0_BASE_ADDR     32'hA000_0000
`define UART0_OFFSET        32'h0000_0FFF