`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Sree Sankar E.
// Create Date: 06.12.2020 11:31:51
// Design Name: RISC V 32I
// Project Name: RISC V Core
// Revision: 1.0
//////////////////////////////////////////////////////////////////////////////////


module top(input i_clk,i_rst);

    risc_core RV32I_core(.i_clk(i_clk),.i_rst(i_rst));

endmodule
