module machine_reg();

endmodule