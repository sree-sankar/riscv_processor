`timescale 1ns / 1ps
//----------------------+-------------------------------------------------------
// Filename             | uart_ctrl.sv
// File created on      | 06/19/2022 18:26:12
// Created by           | Sree Sankar E
//                      |
//                      |
//                      |
//----------------------+-------------------------------------------------------
//
//------------------------------------------------------------------------------
// System Register
//------------------------------------------------------------------------------
module tb_top();

    logic    clk_i    ; // System Clock
    logic    resetn_i ; // Synchronous Active Low System Reset
    // UART
    logic    uart_rx_i;
    logic    uart_tx_o;

//------------------------------------------------------------------------------
// DUT
//------------------------------------------------------------------------------

    top dut(.*);

//------------------------------------------------------------------------------
// DUT
//------------------------------------------------------------------------------

    // Clock
    always #5 clk_i = ~clk_i;

    initial
        begin
        clk_i    <= 'h0;
        resetn_i <= 'h0;
        #20
        resetn_i <= 'h1;
        end

endmodule