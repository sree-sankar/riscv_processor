module mmu (
    ports
);
    
endmodule