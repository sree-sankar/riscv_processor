//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.11.2020 12:07:34
// Design Name: 
// Module Name: define
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//
//
//-----------------Memory Map---------------------------//

`define MEM_MAP_BOOTROM     32'h0000_0000
//`define RESERVED            32'h
`define MEM_MAP_UART0       32'h0000_0000
//`define RESERVED            32'h
`define MEM_MAP_SPI0        32'h0000_0000
`define MEM_MAP_SPI1        32'h0000_0000
//`define RESERVED            32'h
`define MEM_MAP_UART0       32'h0000_0000
//`define RESERVED            32'b
`define MEM_MAP_GPIO0       32'h0000_0000
//`define RESERVED            32'b
`define MEM_MAP_DDR         32'h0000_0000
//`define RESERVED            32'b