module cache_control (
    ports
);
    
endmodule