//----------------------+-------------------------------------------------------
// Filename             | mux2_1_comb.sv
// File created on      | 05.12.2021 08:53:12
// Created by           | Sree Sankar E
//                      |
//                      |
//                      |
//----------------------+-------------------------------------------------------
//
//------------------------------------------------------------------------------
// Adder
//------------------------------------------------------------------------------

module mux2_1_comb#(
    parameter  DW = 32
)(
    input  [DW-1:0]    input0,
    input  [DW-1:0]    input1,
    input              sel   ,
    output [DW-1:0]    result
);

    assign result = (sel) ? input1 : input0;

endmodule