//----------------------+-------------------------------------------------------
// Filename             | shifter.sv
// File created on      | 28.10.2024
// Created by           | Sree Sankar E
//                      |
//                      |
//                      |
//----------------------+-------------------------------------------------------
//
//------------------------------------------------------------------------------
// Shifter
//------------------------------------------------------------------------------

module shifter #(
    parameter DW          = 32 ,
    parameter SHIFT_WIDTH = 5
)(
    input  [   2:0]    opcode_i,
    input  [DW-1:0]    data0_i ,
    input  [DW-1:0]    data1_i ,
    output [DW-1:0]    result_o
);

//------------------------------------------------------------------------------
// Signed
//------------------------------------------------------------------------------

    logic signed [DW-1:0]    data0_signed;
    logic signed [DW-1:0]    sra_res     ;

    assign data0_signed = data0_i;
    assign sra_res      = (data0_signed >>> data1_i[SHIFT_WIDTH-1:0]);

//------------------------------------------------------------------------------
// Output
//------------------------------------------------------------------------------

    assign result_o = (opcode_i[0]) ? (data0_i << data1_i[SHIFT_WIDTH-1:0]) :
                      (opcode_i[1]) ? (data0_i >> data1_i[SHIFT_WIDTH-1:0]) :
                      (opcode_i[2]) ? sra_res : 'h0;

endmodule